module nand_gate (input a, b, output out);

	wire \$n6_0;
	wire \$n5_0;
	wire \$n4_0;

	not (\$n4_0, a);
	not (\$n5_0, b);
	nor (\$n6_0, \$n5_0, \$n4_0);
	not (out, \$n6_0);

endmodule
